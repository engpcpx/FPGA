------------------------------------------------------------------------------
-- exer_02
-- author: Paulo Cezar da Paixao
-- 
------------------------------------------------------------------------------
-- libraries and packages
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
------------------------------------------------------------------------------
-- entity
entity exer_02_view is


   generic(	width :	integer:=8;                             -- memory width
		depth : integer:=8;                             -- memory depth 
		addr  :	integer:=2);                            -- address width

   port (
         clk	 : in  std_logic;				-- clock pulse    
         rst     : in  std_logic;                      	       -- reset memory
         en      : in  std_logic;                               -- enable memory
         d       : in  std_logic;                      	       -- data input
         q_a     : inout  std_logic_vector(7 downto 0);			 -- buffer a
         q_b     : inout  std_logic_vector(7 downto 0); 		    -- buffer b
	      q_c     : inout  std_logic_vector(7 downto 0));        -- buffer c 

end entity;
------------------------------------------------------------------------------
-- architecture
architecture hardware of exer_02_view is



  begin

	process(clk,rst, en)
	begin
	    if rst = '1' then
		 q_a <= (others=>'0'); --x"0"; --x na frende do vetor Ã© HEXA.
		 q_a <= (others=>'0'); --jeito de zerar algo sem saber tamanho.
		 q_c <= (others=>'0');
		 
                 elsif clk'event and clk = '1' then
		       if en = '1' then
			  --jeito 1
			  q_a(0) <= d;
			  q_a(7 downto 1) <= q_a(6 downto 0);
			  --jeito 2: apimentado. igual o jeito 1, mas com uma
			  --constante para o tamanho.
			  q_b(0) <= d;
			  q_b(q_b'high downto 1) <= q_b(q_a'high-1 downto 0);
			  --jeito 3
			  q_c <= q_c(q_c'high-1 downto 0) & d;
			end if;
	      end if;
	end process;
end architecture;