---------------------------------------------------------------------
-- exer 3 - decoder 3to8 using when/else
-- author: Paulo Cezar da Paixao
--
---------------------------------------------------------------------
-- Decodder 3to8 bits
-- using when/else structure
-- 
-- a  b  c    s7 s6 S5 S4 S3 S2	S1 S0
-- 0  0  0    0  0  0  0  0  0  0  1
-- 0  0  1    0  0  0  0  0  0  1  0
-- 0  1  0    0  0  0  0  0  1  0  0
-- 0  1  1    0  0  0  0  1  0  0  0
-- 1  0  0    0  0  0  1  0  0  0  0
-- 1  0  1    0  0  1  0  0  0  0  0 
-- 1  1  0    0  1  0  0  0  0  0  0
-- 1  1  1    1  0  0  0  0  0  0  0

---------------------------------------------------------------------
-- libraries and packages
library ieee;
use ieee.std_logic_1164.all;

---------------------------------------------------------------------
-- entity declaration
entity decoder_3to8_a is 

	port(
		abc :  in  std_logic_vector(2 downto 0);
		s   :  out std_logic_vector(7 downto 0)
	);
		
end decoder_3to8_a;

---------------------------------------------------------------------
-- architecture declaration	
architecture hardware of decoder_3to8_a is

	begin 
		
		s <= 	"00000001" when abc = "000" else
			"00000010" when abc = "001" else
			"00000100" when abc = "010" else
			"00001000" when abc = "011" else
			"00010000" when abc = "100" else
	         	"00100000" when abc = "101" else
			"01000000" when abc = "110" else
			"10000000" when abc = "111";
		
end architecture hardware;